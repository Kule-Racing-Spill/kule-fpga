localparam FRAMEBUFFER_SIZE = 384000;