`ifndef _params_vh
`define _params_vh
localparam FRAMEBUFFER_SIZE = 384000;
`endif