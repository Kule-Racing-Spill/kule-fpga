`timescale 1ns/1ps

module lcd_signals_tb(
    );
endmodule