`timescale 1ns/1ps

module top_tb(
    );
    //vga_signals_tb vga_sig_tb();
    vga_color_tb vga_col_tb();
    framebuffer_tb framebuffer_tb();
endmodule
