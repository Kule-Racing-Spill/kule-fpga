localparam FRAMEBUFFER_SIZE = 192000;